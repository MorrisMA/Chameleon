`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////// 
// Company:         M. A. Morris & Associates
// Engineer:        Michael A. Morris
// 
// Create Date:     12:02:40 10/28/2012 
// Design Name:     WDC W65C02 Microprocessor Re-Implementation
// Module Name:     M65C02_StkPtr.v
// Project Name:    C:\XProjects\ISE10.1i\M65C02A
// Target Devices:  Generic SRAM-based FPGA
// Tool versions:   Xilinx ISE 10.1i SP3
// 
// Description:
//
//  This module implements the functions of the M65C02 stack pointer. The imple-
//  mentation is taken from the M65C02_ALU module so that these functions can be
//  moved to the M65C02_AddrGen module.
//
// Dependencies:    none.
//
// Revision: 
//
//  1.00    13I14   MAM     Implementation pulled from M65C02_ALU. 
//
// Additional Comments: 
//
//  The stack pointer register is a loadable up/down counter. Valid and Rdy are
//  used to generate a local clock enable for the counter. The StkOp input from
//  the microprogram controls the functions implemented. 
//
//  The stack operations supported are: hold, rsvd, ++S, and S--. The stack
//  pointer can only be loaded from the X index register. Similarly, the stack
//  pointer can only be transfered to the X index register. The stack pointer
//  points to an open location on the stack. Thus, push operations write the
//  value at the location pointed to by S, and post-decrements S, S--. Stack 
//  pull operations require the value to be incremented by one, ++S, before
//  that location can be read into OP1 and subsequently written to one of four 
//  registers: P, A, X, or Y.
//
//  The stack pointer control, StkOp, field is generated by the execution
//  engine:
//
//  00  :   Hold;
//  01  :   Rsvd;
//  10  :   S--;
//  11  :   ++S;
//
//  A separate output multiplexer with a built-in incrementer is used to imple-
//  ment the 
//  
//
////////////////////////////////////////////////////////////////////////////////

module M65C02_StkPtr #(
    parameter pStkPtr_Rst = 0
)(
    input   Rst,
    input   Clk,
    
    input   Rdy,
    input   Valid,
    
    input   SelS,
    input   [1:0] Stk_Op,
    input   [7:0] X,
    
    output  reg [7:0] S
);

////////////////////////////////////////////////////////////////////////////////
//
//  Implementation
//

//  Stack Pointer

assign Ld_S = Rdy & (SelS & Valid);
assign CE_S = Rdy & Stk_Op[1];

always @(posedge Clk)
begin
    if(Rst)
        S <= #1 pStkPtr_Rst;
    else if(Ld_S)
        S <= #1 X;                          // TXS
    else if(CE_S)
        S <= #1 ((Stk_Op[0]) ? (S + 1)      // Pop
                             : (S - 1));    // Push
end

endmodule
